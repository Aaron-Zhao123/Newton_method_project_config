library verilog;
use verilog.vl_types.all;
entity Newton_method is
    port(
        x_value         : in     vl_logic_vector(1 downto 0);
        operand_two     : in     vl_logic_vector(1 downto 0);
        subtrahend_one  : in     vl_logic_vector(1 downto 0);
        minuend_one     : in     vl_logic_vector(1 downto 0);
        numerator_one   : in     vl_logic_vector(1 downto 0);
        divisor_one     : in     vl_logic_vector(1 downto 0);
        subtrahend_two  : in     vl_logic_vector(1 downto 0);
        minuend_two     : in     vl_logic_vector(1 downto 0);
        mul_three       : in     vl_logic_vector(1 downto 0);
        subtrahend_three: in     vl_logic_vector(1 downto 0);
        minuend_three   : in     vl_logic_vector(1 downto 0);
        mul_four        : in     vl_logic_vector(1 downto 0);
        operand_four    : in     vl_logic_vector(1 downto 0);
        numerator_two   : in     vl_logic_vector(1 downto 0);
        divisor_two     : in     vl_logic_vector(1 downto 0);
        subtrahend_four : in     vl_logic_vector(1 downto 0);
        minuend_four    : in     vl_logic_vector(1 downto 0);
        clk             : in     vl_logic;
        product_one     : out    vl_logic_vector(1 downto 0);
        product_two     : out    vl_logic_vector(1 downto 0);
        diff_one        : out    vl_logic_vector(1 downto 0);
        quotient_one    : out    vl_logic_vector(1 downto 0);
        diff_two        : out    vl_logic_vector(1 downto 0);
        product_three   : out    vl_logic_vector(1 downto 0);
        diff_three      : out    vl_logic_vector(1 downto 0);
        product_four    : out    vl_logic_vector(1 downto 0);
        quotient_two    : out    vl_logic_vector(1 downto 0);
        diff_four       : out    vl_logic_vector(1 downto 0);
        In_vd_mul_one   : in     vl_logic;
        Out_rd_mul_one  : in     vl_logic;
        In_rd_mul_one   : out    vl_logic;
        Out_vd_mul_one  : out    vl_logic;
        In_vd_sub_one   : in     vl_logic;
        Out_rd_sub_one  : in     vl_logic;
        In_rd_sub_one   : out    vl_logic;
        Out_vd_sub_one  : out    vl_logic;
        In_vd_mul_two   : in     vl_logic;
        Out_rd_mul_two  : in     vl_logic;
        In_rd_mul_two   : out    vl_logic;
        Out_vd_mul_two  : out    vl_logic;
        In_vd_div_one   : in     vl_logic;
        Out_rd_div_one  : in     vl_logic;
        In_rd_div_one   : out    vl_logic;
        Out_vd_div_one  : out    vl_logic;
        In_vd_sub_two   : in     vl_logic;
        Out_rd_sub_two  : in     vl_logic;
        In_rd_sub_two   : out    vl_logic;
        Out_vd_sub_two  : out    vl_logic;
        In_vd_mul_three : in     vl_logic;
        Out_rd_mul_three: in     vl_logic;
        In_rd_mul_three : out    vl_logic;
        Out_vd_mul_three: out    vl_logic;
        In_vd_sub_three : in     vl_logic;
        Out_rd_sub_three: in     vl_logic;
        In_rd_sub_three : out    vl_logic;
        Out_vd_sub_three: out    vl_logic;
        In_vd_mul_four  : in     vl_logic;
        Out_rd_mul_four : in     vl_logic;
        In_rd_mul_four  : out    vl_logic;
        Out_vd_mul_four : out    vl_logic;
        In_vd_div_two   : in     vl_logic;
        Out_rd_div_two  : in     vl_logic;
        In_rd_div_two   : out    vl_logic;
        Out_vd_div_two  : out    vl_logic;
        In_vd_sub_four  : in     vl_logic;
        Out_rd_sub_four : in     vl_logic;
        In_rd_sub_four  : out    vl_logic;
        Out_vd_sub_four : out    vl_logic
    );
end Newton_method;
