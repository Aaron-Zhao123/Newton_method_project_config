library verilog;
use verilog.vl_types.all;
entity testbench_test_handshake is
end testbench_test_handshake;
